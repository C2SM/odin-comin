netcdf station_input {
dimensions:
	obs = unlimited ;
	nchar = 20 ;
variables:
  double stime(obs) ;
    stime:units = "days since 1970-01-01 00:00:00" ;
    stime:long_name = "start time of observation interval; UTC" ;
    stime:calendar = "proleptic_gregorian" ;
  double etime(obs) ;
    etime:units = "days since 1970-01-01 00:00:00" ;
    etime:long_name = "end time of observation interval; UTC" ;
    etime:calendar = "proleptic_gregorian" ;
  float longitude(obs) ;
    longitude:units = "degrees_east";
    longitude:standard_name = "longitude";
    longitude:_FillValue = 1.0e+20f;
  float latitude(obs) ;
    latitude:units = "degrees_north";
    latitude:standard_name = "latitude";
    latitude:_FillValue = 1.0e+20f;
  float elevation(obs) ;
    elevation:units = "m" ;
    elevation:long_name = "surface elevation above sea level" ;
    elevation:_FillValue = 1.0e+20f;
  float sampling_height(obs) ;
    sampling_height:units = "m" ;
    sampling_height:long_name = "sampling height above surface" ;
    sampling_height:_FillValue = 1.0e+20f;
  float sampling_strategy(obs) ;
    sampling_strategy:units = "1" ;
    sampling_strategy:long_name = "sampling strategy flag" ;
    sampling_strategy:comment = "1=low ; 2=mountain ; 3=flight" ;
  char site_name(obs,nchar) ;
    site_name:long_name = "station name or ID" ;

// global attributes:
		:Conventions = "CF-1.8" ;
		:title = "Station input file for ICON ComIn interface XYZ" ;
		:institution = "Empa" ;
		:source = "ICON ComIn interface XYZ" ;
		:version = "1.0" ;
		:author = "Zeno Hug" ;
		:transport_model = "ICON" ;
		:transport_model_version = "" ;
		:experiment = "" ;
		:project = "" ;
		:references = "" ;
		:comment = "" ;
		:license = "CC-BY-4.0" ;
		:history = "" ;
}
